-------------------------------------------------------------------------------
--
-- Title       : sixtyfourbit_module
-- Design      : ALU
-- Author      : riczhang
-- Company     : Stony Brook University
--
-------------------------------------------------------------------------------
--
-- File        : c:\My_Designs\ESE345_PROJECT\ALU\src\sixtyfourbit_module.vhd
-- Generated   : Mon Nov 21 11:00:17 2016
-- From        : interface description file
-- By          : Itf2Vhdl ver. 1.22
--
-------------------------------------------------------------------------------
--
-- Description : 
--
-------------------------------------------------------------------------------

--{{ Section below this comment is automatically maintained
--   and may be overwritten
--{entity {sixtyfourbit_module} architecture {structural}}

library IEEE;
use IEEE.STD_LOGIC_1164.all;

entity sixtyfourbit_module is
end sixtyfourbit_module;

--}} End of automatically maintained section

architecture structural of sixtyfourbit_module is
begin

	 -- enter your statements here --

end structural;
